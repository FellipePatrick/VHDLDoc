library verilog;
use verilog.vl_types.all;
entity teste_vlg_check_tst is
    port(
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end teste_vlg_check_tst;
