library verilog;
use verilog.vl_types.all;
entity teste is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        M1              : out    vl_logic;
        M2              : out    vl_logic;
        M3              : out    vl_logic;
        M4              : out    vl_logic
    );
end teste;
