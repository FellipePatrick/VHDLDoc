library verilog;
use verilog.vl_types.all;
entity teste is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        y               : out    vl_logic
    );
end teste;
